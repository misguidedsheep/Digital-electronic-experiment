library verilog;
use verilog.vl_types.all;
entity DataDistributor_vlg_vec_tst is
end DataDistributor_vlg_vec_tst;
