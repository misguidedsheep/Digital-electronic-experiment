library verilog;
use verilog.vl_types.all;
entity count_vlg_vec_tst is
end count_vlg_vec_tst;
