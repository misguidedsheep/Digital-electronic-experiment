library verilog;
use verilog.vl_types.all;
entity selection2to1_vlg_vec_tst is
end selection2to1_vlg_vec_tst;
