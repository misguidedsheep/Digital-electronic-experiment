library verilog;
use verilog.vl_types.all;
entity lab1 is
    port(
        o3              : out    vl_logic;
        e               : in     vl_logic;
        o2              : out    vl_logic;
        d               : in     vl_logic;
        c               : in     vl_logic;
        o1              : out    vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic
    );
end lab1;
